// Copyright 2019 Politecnico di Torino.
// Copyright and related rights are licensed under the Solderpad Hardware
// License, Version 2.0 (the "License"); you may not use this file except in
// compliance with the License.  You may obtain a copy of the License at
// http://solderpad.org/licenses/SHL-2.0. Unless required by applicable law
// or agreed to in writing, software, hardware and materials distributed under
// this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
// CONDITIONS OF ANY KIND, either express or implied. See the License for the
// specific language governing permissions and limitations under the License.
//
// File: util.svh
// Author: Matteo Perotti
// Date: 02/09/2019

`ifndef UTIL_SVH_
`define UTIL_SVH_

// binary multipliers for Bytes
`define B   *1
`define KiB *1024`B
`define MiB *1024`KiB
`define GiB *1024`MiB
`define TiB *1024`GiB

`endif /* UTIL_SVH_ */